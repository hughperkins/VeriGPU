parameter mem_simulated_delay = 128;
parameter memory_size = 5;
