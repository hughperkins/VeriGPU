/*
Max propagation delay: 70.2 nand units
Area:                  296.0 nand units
*/
module add(input [31:0] a, input [31:0] b, output [31:0] out);
    assign out = a + b;
endmodule
