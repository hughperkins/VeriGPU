parameter width = 32;
