// for use with GLS

parameter mem_simulated_delay = 128;
