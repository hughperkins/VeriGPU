parameter bits_per_cycle = 1;
