// represents a computer, i.e. the combination of processor (proc) and
// memory controller (mem)
module comp(
    input clk,
    input rst,

    input [31:0] oob_wr_addr,
    input [31:0] oob_wr_data,
    input oob_wen,

    output mem_d_req, mem_wr_req,
    output mem_busy,
    output mem_ack,

    output [31:0] out,
    output [6:0] op,
    output [4:0] rd,
    output [6:0] imm1,
    output [31:0] x1,
    output [31:0] pc,
    output [4:0] state,
    output halt,
    output outen
);
    reg [31:0] mem_addr;
    reg [31:0] mem_rd_data, mem_wr_data;

    mem_delayed mem1(
        .clk(clk),

        .addr(mem_addr),
        .wr_req(mem_wr_req), .rd_req(mem_rd_req),
        .rd_data(mem_rd_data), .wr_data(mem_wr_data),
        .busy(mem_busy), .ack(mem_ack),

        .oob_wr_addr(oob_wr_addr), .oob_wr_data(oob_wr_data),
        .oob_wen(oob_wen)
    );

    proc proc1(
        .rst(rst), .clk(clk), .out(out), .op(op), .imm1(imm1), .pc(pc),
        .rd(rd),
        .x1(x1),
        .state(state), .outen(outen), .halt(halt),

        .mem_addr(mem_addr),
        .mem_rd_data(mem_rd_data), .mem_wr_data(mem_wr_data),
        .mem_ack(mem_ack), .mem_busy(mem_busy),
        .mem_rd_req(mem_rd_req), .mem_wr_req(mem_wr_req)
        //.mem_we(mem_we)
    );

endmodule
