/*
use pipeline for int_div, but test writin back to a registry file

required parameters:
- data_width: how many bits in the input and output ints
- num_regs: how many registers there are in the registry file

protocol:
- client wants to divide a by b; and put quotient into register r_quot_sel,
  and modulus into r_mod_sel
- client sets these lines to desired values, and sets req to 1, waits for clock tick
- after clock tick, client sets req to 0
- module takes over
- each clock tick works way through the division
- once done, writes the results to the registers, i.e. quotient then modulus
     - if a register selector is 0, it is ignored,
     - otherwise, for each register, one at a time (different clock ticks):
         - puts selector and data onto rf_wr_sel and rf_wr_data, and sets rf_wr_req; then waits for rf_wr_ack to turn high
         - once rf_wr_ack is high, sets rf_wr_req back to 0
         - if required, continues with modulus, or moves back to IDLE state

$ python toy_proc/timing.py --in-verilog src/int_div_regfile.sv 

Propagation delay is between any pair of combinatorially connected
inputs and outputs, drawn from:
    - module inputs
    - module outputs,
    - flip-flop outputs (treated as inputs), and
    - flip-flop inputs (treated as outputs)

max propagation delay: 44.2 nand units
*/

module int_div_regfile(
    input clk,
    input rst,

    input req,
    output reg busy,

    input [reg_sel_width - 1: 0] r_quot_sel,  // 0 means, dont write (i.e. x0)
    input [reg_sel_width - 1: 0] r_mod_sel,   // 0 means, dont write  (i.e. x0)
    input [data_width - 1:0] a,
    input [data_width - 1:0] b,

    output reg [reg_sel_width - 1:0] rf_wr_sel,
    output reg [data_width - 1:0] rf_wr_data,
    output reg rf_wr_req,
    input rf_wr_ack
);
    parameter data_width = 32;
    parameter num_regs = 32;

    parameter reg_sel_width = $clog2(num_regs);
    parameter pos_width = $clog2(data_width);
    parameter data_width_minus_1 = data_width - 1;

    typedef enum bit[1:0] {
        IDLE,
        CALC,
        WRITING_QUOTIENT,
        WRITING_MODULUS
    } e_state;

    reg [1:0] state;
    reg [pos_width - 1:0] pos;
    reg [data_width - 1:0] quotient;
    reg [data_width - 1:0] remainder;
    reg [data_width - 1: 0] a_remaining;

    reg [1:0] next_state;
    reg [pos_width -1:0] next_pos;
    reg [data_width -1:0] next_quotient;
    reg [data_width -1:0] next_a_remaining;

    reg [reg_sel_width - 1:0] next_rf_wr_sel;
    reg [data_width - 1:0] next_rf_wr_data;
    reg next_rf_wr_req;
    reg next_busy;

    // reg next_ack;

    always @(*) begin
    // always @(state, pos, req, rf_wr_ack) begin
        reg [2 * data_width - 1: 0] shiftedb;

        // rf_wr_req = 0;
        next_state = state;
        next_pos = pos;
        // busy = 0;
        next_quotient = quotient;
        next_a_remaining = a_remaining;
        next_busy = 0;
        // next_ack = 0;

        next_rf_wr_req = 0;
        next_rf_wr_sel = '0;
        next_rf_wr_data = '0;

        shiftedb = {{data_width{1'b0}}, b} << pos;

        $display("div comb req=%0d state=%0d pos=%0d rf_wr_ack=%0d", req, state, pos, rf_wr_ack);
        // $strobe("state %0d req=%0b", state, req);
        case(state)
            IDLE: begin
                if(req) begin
                    $display("div unit got req");
                    next_pos = data_width_minus_1[pos_width - 1:0];
                    next_quotient = '0;
                    next_a_remaining = a;
                    next_busy = 1;
                    next_state = CALC;
                end
            end
            CALC: begin
                next_busy = 1;
                if (shiftedb < {{data_width{1'b0}}, next_a_remaining}) begin
                    next_a_remaining = next_a_remaining - shiftedb[data_width - 1 :0];
                    next_quotient[pos] = 1;
                end
                if (pos == 0) begin
                    if(r_quot_sel != 0) begin
                        next_rf_wr_req = 1;
                        next_rf_wr_sel = r_quot_sel;
                        next_rf_wr_data = next_quotient;
                        next_state = WRITING_QUOTIENT;
                        $display("div. wrote quotient");
                    end else if(r_mod_sel != 0) begin
                        next_rf_wr_req = 1;
                        next_rf_wr_sel = r_mod_sel;
                        next_rf_wr_data = next_a_remaining;
                        next_state = WRITING_MODULUS;
                    end else begin
                        next_state = IDLE;  // this should never normally happen :), but it's a possible input
                    end
                end else begin
                    next_pos = pos - 1;
                end
            end
            WRITING_QUOTIENT: begin
                if(rf_wr_ack) begin
                    $display("div got ack, maybe write modulus");
                    if(r_mod_sel != 0) begin
                        $display("div write modulus (for next cycle)");
                        next_busy = 1;
                        next_rf_wr_req = 1;
                        next_rf_wr_sel = r_mod_sel;
                        next_rf_wr_data = next_a_remaining;
                        next_state = WRITING_MODULUS;
                    end else begin
                        next_state = IDLE;
                    end
                end else begin
                    $display("div waiting ack");
                    next_busy = 1;
                    next_rf_wr_req = 1;
                    next_rf_wr_sel = r_quot_sel;
                    next_rf_wr_data = next_quotient;
                end
            end
            WRITING_MODULUS: begin
                if(rf_wr_ack) begin
                    next_state = IDLE;
                end else begin
                    next_busy = 1;
                    next_rf_wr_req = 1;
                    next_rf_wr_sel = r_mod_sel;
                    next_rf_wr_data = next_a_remaining;
                end
            end
        endcase
    end

    always @(posedge clk, posedge rst) begin
        // $strobe("always %0d req=%0b rst=%0b", state, req, rst);
        if (rst) begin
            state <= IDLE;
            pos <= 0;
            busy <= 0;

            rf_wr_req <= 0;
            rf_wr_sel <= 0;
            rf_wr_data <= 0;
            busy <= 0;
            // ack <= 0;
        end else begin
            // $display("div clk");
            state <= next_state;
            pos <= next_pos;
            quotient <= next_quotient;
            a_remaining <= next_a_remaining;

            rf_wr_req <= next_rf_wr_req;
            rf_wr_sel <= next_rf_wr_sel;
            rf_wr_data <= next_rf_wr_data;

            busy <= next_busy;
            // ack <= next_ack;
        end
    end
endmodule
