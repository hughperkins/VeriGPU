/*
experiment with various parallel adds
*/
module mul_partial_add(
    input [23:0] a,
    input [23:0] b,
    output reg [47:0] out [4]
);
endmodule
