// test assign with timing.py
module test_assign(input [2:0] a, output [2:0] out);
    assign out = a;
endmodule
