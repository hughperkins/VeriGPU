`define assert_known(VAL) begin end

`define assert(VAL) begin end
